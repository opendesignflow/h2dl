module LongFileModule (

    input clk,
    input res_n,
    
    input wire a,
    
    input wire [7:0] a,
    
    output wire a, 
    
    output reg b,
    
    output reg [7:0] c
);


    // A
    //---------
    
    // B
    //-------------



endmodule